module segment_show(input clock,input reset,input [11:0]data_show,
input [2:0]byte_status,output [3:0]bytee,output[6:0]segment,input [3:0]segment_byte_control);

endmodule
